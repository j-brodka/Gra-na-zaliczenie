0 0 30 1 3 10
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1
1

0
0
0
0

